`timescale 1ns/1ps

//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date:    10:58:01 10/10/2011
// Design Name:
// Module Name:    alu_top
// Project Name:
// Target Devices:
// Tool versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////

module alu_top(
               src1,       //1 bit source 1 (input)
               src2,       //1 bit source 2 (input)
               less,       //1 bit less     (input)
               A_invert,   //1 bit A_invert (input)
               B_invert,   //1 bit B_invert (input)
               cin,        //1 bit carry in (input)
               operation,  //operation      (input)
               result,     //1 bit result   (output)
               cout,       //1 bit carry out(output)
               );

input         src1;
input         src2;
input         less;
input         A_invert;
input         B_invert;
input         cin;
input [2-1:0] operation;

output        result;
output        cout;

reg           result;

always@( * )
begin
    if ( A_invert ) begin
        A = ~src1;
    end
    else begin
        A = src1;
    end

    if ( B_invert ) begin
        B = ~src2;
    end
    else begin
        B = src2;
    end

    case(operation)
    2'd0:  begin
        result <= A & B;
    end

    2'd1:  begin
        result <= A | B;
    end

    2'd2:  begin
        result <= (A&B) | (cin&B) | (cin&A);
    end

    2'd3:  begin

    end
    endcase
end

endmodule
